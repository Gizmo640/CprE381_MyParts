library IEEE;
use IEEE.std_logic_1164.all;

entity Decoder_5t32 is
	port(
		Enable_Signal: in STD_LOGIC;
		Input_In: in std_logic_vector(4 downto 0);
		Output_Out: out std_logic_vector(31 downto 0));
end Decoder_5t32;

architecture Design of Decoder_5t32 is
begin
	Output_Out <=
		"00000000000000000000000000000000" when (Enable_Signal = '0') else
		"00000000000000000000000000000001" when (Input_In = "00000") else
		"00000000000000000000000000000010" when (Input_In = "00001") else
		"00000000000000000000000000000100" when (Input_In = "00010") else
		"00000000000000000000000000001000" when (Input_In = "00011") else
		"00000000000000000000000000010000" when (Input_In = "00100") else
		"00000000000000000000000000100000" when (Input_In = "00101") else
		"00000000000000000000000001000000" when (Input_In = "00110") else
		"00000000000000000000000010000000" when (Input_In = "00111") else
		"00000000000000000000000100000000" when (Input_In = "01000") else
		"00000000000000000000001000000000" when (Input_In = "01001") else
		"00000000000000000000010000000000" when (Input_In = "01010") else
		"00000000000000000000100000000000" when (Input_In = "01011") else
		"00000000000000000001000000000000" when (Input_In = "01100") else
		"00000000000000000010000000000000" when (Input_In = "01101") else
		"00000000000000000100000000000000" when (Input_In = "01110") else
		"00000000000000001000000000000000" when (Input_In = "01111") else
		"00000000000000010000000000000000" when (Input_In = "10000") else
		"00000000000000100000000000000000" when (Input_In = "10001") else
		"00000000000001000000000000000000" when (Input_In = "10010") else
		"00000000000010000000000000000000" when (Input_In = "10011") else
		"00000000000100000000000000000000" when (Input_In = "10100") else
		"00000000001000000000000000000000" when (Input_In = "10101") else
		"00000000010000000000000000000000" when (Input_In = "10110") else
		"00000000100000000000000000000000" when (Input_In = "10111") else
		"00000001000000000000000000000000" when (Input_In = "11000") else
		"00000010000000000000000000000000" when (Input_In = "11001") else
		"00000100000000000000000000000000" when (Input_In = "11010") else
		"00001000000000000000000000000000" when (Input_In = "11011") else
		"00010000000000000000000000000000" when (Input_In = "11100") else
		"00100000000000000000000000000000" when (Input_In = "11101") else
		"01000000000000000000000000000000" when (Input_In = "11110") else
		"10000000000000000000000000000000" when (Input_In = "11111") else
		(31 downto 0 => '0');
end Design;