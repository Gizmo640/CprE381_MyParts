library IEEE;
use IEEE.std_logic_1164.all;

package MyPackage is
	type STD_LOGIC_ARRAY is array (natural range <>) of STD_LOGIC_VECTOR;

end package MyPackage;
